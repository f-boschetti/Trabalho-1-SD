-- teste de commit

--###########################
--#   VER COM O PROFESSOR   #
--###########################


--N�o entendi como implementar o multiplicador no projeto
--Provavelmente vai ser preciso colocar todos os projetos em um arquivo s� pois n�o sei como funciona
-- o sistema para importar "component" em VHDL, talvez ele considere tudo do mesmo diretorio, porem n�o encontrei nada
--na internet

--mas uma possibilidade � copiar todos os codigos em um s� 


--primeiro
	--fazer a descri��o completa de todos os componentes "menores" com entity e architecture normal,
	--exatamente igual aos projetos originais

--segundo
	-- fazer o projeto "maior" e declarar na architecture os componentes e seus port maps
	-- (isso antes dos sinais e do begin da architecture)
	
--terceiro 
	--fazer o port map dos sinais depois do begin da architecture
	
	
	
-- OUTRA OP��O � tambem usar como function, porem eu nao pesquisei como usar ainda